magic
tech scmos
timestamp 1699601116
<< metal1 >>
rect 89 113 150 122
rect 131 94 140 113
rect 81 62 113 67
rect 108 57 113 62
rect 108 53 124 57
rect 168 52 194 57
rect 15 22 28 30
rect 56 24 59 29
rect -6 13 1 20
rect 128 13 134 19
rect -6 7 155 13
use not  not_0
timestamp 1698904140
transform 1 0 133 0 1 28
box -15 -9 48 66
use nand  nand_0
timestamp 1698951989
transform 1 0 34 0 1 19
box -48 1 68 103
<< labels >>
rlabel metal1 188 54 189 55 1 out
rlabel metal1 19 25 20 27 1 a
rlabel metal1 57 25 58 27 1 b
rlabel metal1 128 115 132 117 1 vdd
rlabel metal1 73 8 76 10 1 gnd
<< end >>
