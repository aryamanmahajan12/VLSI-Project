* SPICE3 file created from fand.ext - technology: scmos



.include TSMC_180nm.txt

.option scale=0.09u


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'



Vin1 in1 gnd DC 1.8

Vin2 in2 gnd DC 1.8

Vin3 in3 gnd DC 1.8

Vin4 in4 gnd DC 1.8

Vin5 in5 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 80ns)

















.option scale=0.09u

M1000 a_n24_n100# in2 a_n74_n100# Gnd CMOSN w=29 l=9
+  ad=1131 pd=136 as=1189 ps=140
M1001 out in1 vdd w_n133_43# CMOSP w=28 l=9
+  ad=3108 pd=390 as=3806 ps=498
M1002 out in5 vdd w_n133_43# CMOSP w=28 l=9
+  ad=0 pd=0 as=0 ps=0
M1003 a_70_n100# in4 a_24_n100# Gnd CMOSN w=29 l=9
+  ad=957 pd=124 as=1073 ps=132
M1004 vdd in2 out w_n133_43# CMOSP w=28 l=9
+  ad=0 pd=0 as=0 ps=0
M1005 a_n74_n100# in1 gnd Gnd CMOSN w=29 l=9
+  ad=0 pd=0 as=1959 ps=250
M1006 out in5 a_70_n100# Gnd CMOSN w=29 l=9
+  ad=986 pd=126 as=0 ps=0
M1007 out1 out vdd w_194_44# CMOSP w=22 l=30
+  ad=902 pd=126 as=0 ps=0
M1008 a_24_n100# in3 a_n24_n100# Gnd CMOSN w=29 l=9
+  ad=0 pd=0 as=0 ps=0
M1009 out1 out gnd Gnd CMOSN w=31 l=30
+  ad=2573 pd=228 as=0 ps=0
M1010 out in3 vdd w_n133_43# CMOSP w=28 l=9
+  ad=0 pd=0 as=0 ps=0
M1011 vdd in4 out w_n133_43# CMOSP w=28 l=9
+  ad=0 pd=0 as=0 ps=0
C0 w_n133_43# vdd 0.15fF
C1 w_194_44# out 0.68fF
C2 w_n133_43# in2 0.22fF
C3 out in5 0.41fF
C4 w_n133_43# in4 0.22fF
C5 w_194_44# vdd 0.12fF
C6 w_n133_43# in3 0.22fF
C7 in2 out 0.41fF
C8 w_194_44# out1 0.12fF
C9 out in4 0.41fF
C10 w_n133_43# in5 0.22fF
C11 w_n133_43# in1 0.22fF
C12 w_n133_43# out 0.19fF
C13 in3 out 0.41fF
C14 gnd Gnd 3.78fF
C15 out1 Gnd 0.94fF
C16 out Gnd 7.84fF
C17 vdd Gnd 3.40fF
C18 in5 Gnd 1.55fF
C19 in4 Gnd 1.55fF
C20 in3 Gnd 1.55fF
C21 in2 Gnd 1.55fF
C22 in1 Gnd 0.09fF
C23 w_194_44# Gnd 5.23fF
C24 w_n133_43# Gnd 12.77fF


*replace text


.tran 1n 800n

.control

run
set color0 = rgb:f/f/e
set color1 = black

plot v(in1) v(in2)+2 v(in3)+4 v(in4)+6 v(in5)+8 v(out1)+10
quit

.end
.endc