magic
tech scmos
timestamp 1699989160
<< metal1 >>
rect 139 965 163 970
rect 139 946 1435 965
rect 1820 951 2724 968
rect 139 245 163 946
rect 2712 866 2724 951
rect 1854 822 2688 828
rect 2665 809 2688 822
rect 2812 811 2826 818
rect 2665 797 2793 809
rect 1460 728 1479 745
rect 1511 730 1527 746
rect 1557 731 1575 745
rect 1605 732 1620 745
rect 1651 734 1726 746
rect 808 713 909 714
rect 808 689 814 713
rect 850 689 1439 713
rect 2740 704 2761 749
rect 1879 690 2773 704
rect 908 688 1439 689
rect -139 188 0 197
rect 680 192 912 204
rect 1592 190 1864 200
rect -29 -124 -25 188
rect 2544 175 2827 185
rect 59 139 67 140
rect 103 133 105 140
rect 970 112 978 113
rect 1929 100 1930 107
rect 2885 96 2893 97
rect 2921 96 2929 97
rect 680 -2 692 1
rect 680 -18 735 -2
rect 756 -18 814 -2
rect 850 -18 1317 -2
rect 1605 -26 2269 -13
rect 2557 -32 3232 -24
rect -29 -138 170 -124
rect -29 -148 -25 -138
rect 164 -173 170 -138
rect 225 -179 1085 -174
rect 1080 -184 1088 -179
rect 1525 -181 1970 -180
rect 1149 -186 1970 -181
rect 2030 -184 3067 -178
rect 2036 -187 3067 -184
rect 2945 -201 2948 -187
rect 161 -216 170 -210
rect 214 -215 225 -210
rect 1138 -222 1161 -217
rect 2019 -221 2050 -216
rect 227 -248 724 -242
rect 756 -244 853 -242
rect 756 -248 1085 -244
rect 853 -249 1085 -248
rect 1075 -255 1089 -249
rect -32 -270 225 -259
rect 1156 -267 1161 -222
rect 1313 -255 1970 -249
rect 2038 -260 2047 -221
rect 2995 -243 3032 -238
rect 2133 -247 2914 -246
rect 2152 -253 2914 -247
rect 1939 -266 2047 -260
rect 990 -268 1161 -267
rect -32 -429 -21 -270
rect 982 -273 1161 -268
rect 982 -274 1156 -273
rect 982 -275 1075 -274
rect 983 -343 990 -275
rect 946 -356 990 -343
rect -30 -643 -21 -429
rect 451 -499 563 -488
rect 59 -597 69 -580
rect 102 -598 125 -579
rect 102 -608 110 -598
rect 121 -608 125 -598
rect 159 -596 168 -580
rect 206 -597 216 -580
rect 206 -605 208 -597
rect 214 -605 216 -597
rect 248 -596 256 -579
rect -30 -654 110 -643
rect 121 -654 126 -643
rect 528 -984 546 -499
rect 949 -589 958 -356
rect 1659 -357 1724 -340
rect 1417 -477 1560 -465
rect 1025 -577 1039 -562
rect 1077 -580 1089 -561
rect 1128 -585 1137 -562
rect 949 -596 951 -589
rect 1174 -580 1183 -562
rect 1217 -573 1280 -561
rect 1174 -590 1176 -580
rect 949 -599 958 -596
rect 1128 -856 1145 -638
rect 1176 -727 1188 -639
rect 526 -2278 546 -984
rect 1525 -1076 1547 -477
rect 1935 -583 1944 -266
rect 2911 -271 2914 -253
rect 2911 -277 2946 -271
rect 2358 -358 2954 -344
rect 2968 -357 3006 -344
rect 2968 -358 3018 -357
rect 2481 -480 2520 -456
rect 2392 -492 2520 -480
rect 2001 -576 2010 -564
rect 2047 -583 2060 -563
rect 2100 -585 2109 -564
rect 2143 -594 2155 -564
rect 2188 -583 2197 -563
rect 2188 -587 2250 -583
rect 2256 -587 2258 -583
rect 2143 -597 2270 -594
rect 2113 -709 2131 -691
rect 2101 -763 2131 -709
rect 2101 -784 2102 -763
rect 815 -1079 1547 -1076
rect 815 -1113 850 -1079
rect 884 -1113 1547 -1079
rect 815 -1114 1525 -1113
rect 2481 -1138 2520 -492
rect 1655 -2096 2263 -2047
rect 1655 -2097 2294 -2096
rect 1705 -2256 1706 -2251
rect 525 -2302 546 -2278
rect 525 -2316 1325 -2302
rect 525 -2343 546 -2316
rect 1357 -2324 1374 -2310
rect 1406 -2324 1422 -2310
rect 1427 -2324 1429 -2310
rect 1452 -2323 1495 -2313
rect 2497 -2440 2520 -1138
rect 2735 -2002 2794 -358
rect 3024 -485 3032 -243
rect 3053 -344 3068 -187
rect 3053 -359 3068 -357
rect 2901 -494 3032 -485
rect 2902 -635 2910 -494
rect 3136 -649 3142 -583
rect 3118 -1245 3144 -649
rect 3117 -1246 3144 -1245
rect 3117 -1841 3143 -1246
rect 2735 -2094 2736 -2002
rect 2793 -2094 2794 -2002
rect 2735 -2095 2794 -2094
rect 3115 -1842 3143 -1841
rect 1427 -2465 2520 -2440
rect 3115 -2303 3141 -1842
rect 3140 -2328 3141 -2303
rect 3115 -2493 3141 -2328
<< m2contact >>
rect 1720 951 1725 970
rect 2805 811 2812 818
rect 2863 802 2871 809
rect 1460 722 1479 728
rect 1511 718 1527 730
rect 1557 725 1575 731
rect 1605 725 1620 732
rect 814 689 850 713
rect 731 61 736 66
rect 1639 34 1648 39
rect 2592 28 2600 33
rect 3556 18 3563 23
rect 814 -18 850 -2
rect 225 -215 234 -210
rect 1137 -255 1151 -249
rect 225 -270 234 -259
rect 1292 -255 1313 -249
rect 2016 -253 2032 -248
rect 2133 -253 2152 -247
rect 405 -366 417 -355
rect 110 -608 121 -598
rect 159 -609 168 -596
rect 208 -605 214 -597
rect 248 -608 256 -596
rect 462 -634 476 -619
rect 110 -654 121 -643
rect 1001 -366 1014 -346
rect 1280 -356 1287 -337
rect 1359 -356 1386 -340
rect 1645 -357 1659 -340
rect 1724 -357 1737 -340
rect 1077 -587 1089 -580
rect 951 -596 958 -589
rect 1128 -594 1137 -585
rect 1280 -573 1286 -561
rect 1176 -590 1183 -580
rect 1005 -613 1039 -601
rect 1128 -638 1145 -630
rect 1176 -639 1188 -634
rect 1176 -751 1188 -727
rect 1128 -907 1145 -856
rect 1973 -357 1986 -340
rect 2250 -358 2256 -339
rect 2270 -358 2276 -339
rect 2954 -358 2968 -344
rect 3006 -357 3018 -344
rect 1935 -597 1944 -583
rect 2047 -597 2060 -583
rect 2101 -593 2109 -585
rect 2250 -591 2256 -583
rect 2270 -597 2276 -583
rect 2101 -709 2113 -691
rect 2102 -784 2131 -763
rect 850 -1113 884 -1079
rect 2263 -2096 2294 -2046
rect 1706 -2256 1713 -2251
rect 1374 -2324 1394 -2310
rect 1422 -2324 1427 -2310
rect 1495 -2323 1508 -2313
rect 3053 -357 3068 -344
rect 2954 -521 2968 -513
rect 2999 -619 3011 -611
rect 2902 -643 2910 -635
rect 2736 -2094 2793 -2002
rect 1422 -2465 1427 -2440
rect 3115 -2328 3140 -2303
<< metal2 >>
rect 741 739 752 752
rect 741 729 1427 739
rect 1720 734 1725 951
rect 741 66 752 729
rect 1421 728 1427 729
rect 1421 722 1460 728
rect 1509 718 1511 730
rect 1527 718 1529 730
rect 736 61 749 66
rect 814 -2 850 689
rect 1509 653 1529 718
rect 1557 677 1575 725
rect 1605 717 1620 725
rect 1604 710 1974 717
rect 1557 666 1755 677
rect 1679 653 1695 654
rect 1509 638 1695 653
rect 1679 39 1695 638
rect 1733 424 1755 666
rect 1948 487 1974 710
rect 2805 646 2812 811
rect 2863 809 2871 829
rect 2805 630 3702 646
rect 3578 487 3586 492
rect 1946 459 3586 487
rect 2662 424 2671 439
rect 1734 400 2671 424
rect 1648 34 1722 39
rect 225 -259 234 -215
rect 1151 -255 1292 -249
rect 405 -355 1001 -346
rect 417 -366 1001 -355
rect 1280 -561 1287 -356
rect 1386 -356 1645 -340
rect 1359 -357 1645 -356
rect 1286 -573 1287 -561
rect 1077 -589 1089 -587
rect 958 -596 1089 -589
rect 110 -643 121 -608
rect 149 -609 159 -596
rect 168 -609 173 -596
rect 149 -856 173 -609
rect 208 -727 214 -605
rect 256 -608 258 -596
rect 248 -644 258 -608
rect 985 -613 1005 -601
rect 985 -618 1039 -613
rect 462 -619 724 -618
rect 476 -634 724 -619
rect 756 -632 1039 -618
rect 1128 -630 1145 -594
rect 756 -634 985 -632
rect 1176 -634 1188 -590
rect 1687 -643 1694 34
rect 2662 33 2671 400
rect 2600 28 2675 33
rect 2016 -248 2133 -247
rect 2032 -253 2133 -248
rect 1737 -357 1973 -340
rect 2250 -583 2256 -358
rect 1944 -597 2047 -583
rect 2060 -597 2062 -583
rect 2109 -593 2113 -585
rect 2270 -583 2276 -358
rect 1218 -644 1694 -643
rect 248 -656 1694 -644
rect 248 -665 1219 -656
rect 1687 -659 1694 -656
rect 2101 -691 2113 -593
rect 2661 -727 2671 28
rect 3578 23 3586 459
rect 3563 18 3590 23
rect 3018 -357 3053 -344
rect 2954 -513 2968 -358
rect 2999 -635 3011 -619
rect 2910 -643 3011 -635
rect 208 -751 1176 -727
rect 1188 -744 2671 -727
rect 1188 -751 2661 -744
rect 2102 -856 2132 -784
rect 3570 -856 3589 18
rect -30 -907 1128 -856
rect 1145 -907 3589 -856
rect 3570 -908 3589 -907
rect 850 -2407 883 -1113
rect 2264 -2046 2736 -2003
rect 2294 -2094 2736 -2046
rect 2294 -2096 2792 -2094
rect 2264 -2109 2792 -2096
rect 3697 -2251 3702 630
rect 1713 -2256 3703 -2251
rect 1374 -2335 1394 -2324
rect 1356 -2343 1394 -2335
rect 1519 -2313 3115 -2303
rect 1508 -2323 3115 -2313
rect 849 -2426 883 -2407
rect 850 -2446 883 -2426
rect 1356 -2446 1373 -2343
rect 1422 -2440 1427 -2324
rect 1519 -2328 3115 -2323
rect 850 -2464 1368 -2446
<< m3contact >>
rect 724 -634 756 -618
<< m123contact >>
rect 59 133 67 139
rect 97 133 103 140
rect 970 106 978 112
rect 1007 106 1015 113
rect 1922 100 1929 107
rect 1958 100 1966 107
rect 735 -18 756 -2
rect 155 -216 161 -210
rect 1094 -223 1103 -217
rect 724 -248 756 -242
rect 1025 -585 1039 -577
rect 59 -609 69 -597
rect 1413 -616 1445 -604
rect 2885 90 2893 96
rect 2921 90 2929 96
rect 1975 -222 1984 -216
rect 1995 -576 2001 -564
rect 1976 -616 1998 -604
rect 2397 -619 2417 -603
rect 2951 -244 2961 -238
rect 2963 -613 2976 -602
rect 2964 -628 2972 -622
rect 1260 -2425 1286 -2407
<< metal3 >>
rect 59 -335 67 133
rect 97 -209 103 133
rect 969 106 970 112
rect 735 -110 756 -18
rect 97 -210 161 -209
rect 97 -216 155 -210
rect -8 -343 67 -335
rect -8 -597 -1 -343
rect 59 -344 67 -343
rect 724 -242 756 -110
rect -8 -609 59 -597
rect 69 -609 70 -597
rect 724 -618 756 -248
rect 969 -577 978 106
rect 1007 -217 1015 106
rect 1007 -223 1094 -217
rect 1922 -564 1929 100
rect 1958 -216 1966 100
rect 2885 23 2893 90
rect 1958 -222 1975 -216
rect 1958 -223 1984 -222
rect 1958 -224 1966 -223
rect 1922 -576 1995 -564
rect 969 -585 1025 -577
rect 969 -586 978 -585
rect 2886 -602 2893 23
rect 2921 -238 2929 90
rect 2921 -244 2951 -238
rect 2397 -603 2841 -602
rect 1445 -616 1976 -604
rect 2417 -619 2841 -603
rect 2886 -613 2963 -602
rect 724 -2405 756 -634
rect 2828 -653 2841 -619
rect 2964 -653 2972 -628
rect 2828 -662 2982 -653
rect 724 -2407 1284 -2405
rect 724 -2425 1260 -2407
rect 724 -2428 756 -2425
use or  or_0
timestamp 1699074691
transform 1 0 1374 0 1 -2214
box -131 -212 331 137
use fand  fand_3
timestamp 1699037659
transform 1 0 144 0 1 -478
box -133 -157 351 123
use xnor  xnor_0
timestamp 1699893713
transform 1 0 0 0 1 34
box 0 -34 737 232
use not  not_0
timestamp 1698904140
transform 1 0 179 0 1 -239
box -15 -9 48 66
use fand  fand_1
timestamp 1699037659
transform 1 0 1113 0 1 -460
box -133 -157 351 123
use not  not_1
timestamp 1698904140
transform 1 0 1103 0 1 -246
box -15 -9 48 66
use xnor  xnor_1
timestamp 1699893713
transform 1 0 912 0 1 7
box 0 -34 737 232
use fand  fand_2
timestamp 1699037659
transform 1 0 2085 0 1 -462
box -133 -157 351 123
use not  not_2
timestamp 1698904140
transform 1 0 1984 0 1 -245
box -15 -9 48 66
use xnor  xnor_2
timestamp 1699893713
transform 1 0 1864 0 1 1
box 0 -34 737 232
use and  and_0
timestamp 1699601116
transform 1 0 2948 0 1 -635
box -14 7 194 122
use not  not_3
timestamp 1698904140
transform 1 0 2960 0 1 -267
box -15 -9 48 66
use xnor  xnor_3
timestamp 1699893713
transform 1 0 2827 0 1 -9
box 0 -34 737 232
use fand  fand_0
timestamp 1699037659
transform 1 0 1547 0 1 847
box -133 -157 351 123
use tor  tor_0
timestamp 1699809212
transform 1 0 2802 0 1 800
box -90 -51 158 73
<< labels >>
rlabel metal1 1863 824 1864 825 1 out
rlabel metal1 150 778 153 780 1 vdd
rlabel metal1 922 697 925 699 1 gnd
rlabel metal1 61 135 62 136 1 a0
rlabel metal1 99 135 100 136 1 b0
rlabel metal1 973 108 974 109 1 a1
rlabel metal1 1010 108 1011 109 1 b1
rlabel metal1 1924 102 1925 103 1 a2
rlabel metal1 1961 102 1962 103 1 b2
rlabel metal1 2887 92 2888 93 1 a3
rlabel metal1 2923 93 2924 94 1 b3
rlabel m2contact 1709 -2254 1710 -2253 1 s1
rlabel metal1 1111 -1097 1113 -1095 1 d1
rlabel metal1 2497 -1086 2499 -1083 1 d2
rlabel metal1 3132 -1038 3134 -1035 1 d3
rlabel metal2 2864 817 2865 818 1 s2
<< end >>
