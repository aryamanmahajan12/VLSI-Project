magic
tech scmos
timestamp 1698904140
<< nwell >>
rect -15 38 46 59
<< ntransistor >>
rect 14 8 18 14
<< ptransistor >>
rect 14 45 18 52
<< ndiffusion >>
rect 8 8 14 14
rect 18 8 23 14
<< pdiffusion >>
rect 8 45 14 52
rect 18 45 23 52
<< ndcontact >>
rect 4 8 8 14
rect 23 8 28 14
<< pdcontact >>
rect 4 45 8 52
rect 23 45 28 52
<< polysilicon >>
rect 14 52 18 56
rect 14 29 18 45
rect 7 23 18 29
rect 14 14 18 23
rect 14 5 18 8
<< polycontact >>
rect 2 23 7 29
<< metal1 >>
rect -15 59 46 66
rect 4 52 8 59
rect 23 29 28 45
rect -9 23 2 29
rect 23 24 35 29
rect 23 14 28 24
rect 4 -3 8 8
rect -14 -9 48 -3
<< labels >>
rlabel metal1 14 61 16 62 5 vdd
rlabel metal1 32 27 34 28 1 out
rlabel metal1 31 -7 33 -6 1 gnd
rlabel metal1 -5 25 -3 27 1 in
<< end >>
