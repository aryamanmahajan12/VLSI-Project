* SPICE3 file created from not.ext - technology: scmos
.include TSMC_180nm.txt

.option scale=0.09u


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'

Vin in gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)

M1000 out in vdd vdd CMOSP w=7 l=4
+  ad=70 pd=34 as=70 ps=34
M1001 out in gnd Gnd CMOSN w=6 l=4
+  ad=60 pd=32 as=60 ps=32

C0 vdd out 0.04fF
C1 vdd in 0.11fF
C2 out vdd 0.03fF
C3 vdd vdd 0.09fF
C4 gnd Gnd 0.18fF
C5 out Gnd 0.12fF
C6 vdd Gnd 0.08fF
C7 in Gnd 0.38fF
C8 vdd Gnd 1.29fF



.measure tran trise 
+ TRIG v(in) VAL = 'SUPPLY/2' RISE =1
+ TARG v(out) VAL = 'SUPPLY/2' RISE =1 

.measure tran tfall 
+ TRIG v(in) VAL = 'SUPPLY/2' FALL =1 
+ TARG v(out) VAL = 'SUPPLY/2' FALL =1



.measure tran tpd param = '(trise + tfall)/2' goal = 0
        

.tran 1n 800n

.control

run
set color0 = rgb:f/f/e
set color1 = black

plot v(in) v(out)+2


quit

.end
.endc