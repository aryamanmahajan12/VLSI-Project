magic
tech scmos
timestamp 1701531022
<< metal1 >>
rect 12306 6807 13117 6822
rect 11643 6770 11684 6773
rect 12308 6771 12312 6776
rect 11643 6766 12062 6770
rect 11643 6751 11684 6766
rect 12055 6758 12062 6766
rect 12055 6752 12174 6758
rect 11980 6742 12141 6749
rect 11980 6717 11994 6742
rect 11601 6704 11997 6717
rect 13048 5657 13117 6807
rect 12511 5638 13117 5657
rect 12566 5481 12570 5486
rect 8601 5254 8634 5255
rect 8374 5245 8634 5254
rect 1244 4604 1385 4610
rect 1244 4165 1268 4604
rect 1580 4543 8699 4548
rect 1351 4498 1366 4503
rect 1375 4498 1380 4503
rect 3013 4023 3021 4029
rect 4065 4026 4069 4031
rect 8673 3732 8685 4543
rect 13048 4181 13117 5638
rect 12665 4178 13117 4181
rect 12664 4158 13117 4178
rect 12719 4001 12723 4006
rect 12156 3937 12303 3947
rect 12147 3926 12303 3937
rect 12147 3732 12156 3926
rect 8673 3716 12157 3732
rect 8123 3637 8124 3654
rect 8132 3637 12381 3654
rect 4612 3394 5351 3397
rect 5756 3394 7662 3397
rect 13048 3395 13117 4158
rect 13000 3394 13117 3395
rect 4612 3388 13117 3394
rect 7656 3387 13117 3388
rect 785 3208 792 3209
rect -3242 2804 -3241 2809
rect -9782 2789 -9781 2794
rect -2150 2593 -1864 2601
rect -2190 2557 -2185 2562
rect -10356 2291 -10350 2300
rect -10797 1906 -10764 1909
rect -10765 1876 -10764 1906
rect -10797 1281 -10764 1876
rect -6598 1763 -6560 1764
rect -8055 1711 -8051 1717
rect -10378 1689 -10374 1695
rect -10772 1235 -10764 1281
rect -10377 992 -10372 1660
rect -8893 1324 -8871 1649
rect -8059 1192 -8053 1683
rect -6598 1356 -6560 1729
rect -5919 1725 -5915 1731
rect -3824 1719 -3820 1725
rect -5926 1424 -5919 1700
rect -4476 1579 -4471 1667
rect -3824 1583 -3817 1687
rect -3824 1582 -3154 1583
rect -3824 1574 -3149 1582
rect -3153 1481 -3149 1574
rect -3419 1424 -3413 1436
rect -5936 1418 -3413 1424
rect -3686 1192 -3681 1202
rect -8060 1174 -3681 1192
rect -3989 992 -3984 1016
rect -10377 988 -3984 992
rect -10376 969 -3984 988
rect -3989 595 -3984 969
rect -3686 598 -3681 1174
rect -3419 595 -3413 1418
rect -3414 587 -3413 595
rect -3152 509 -3148 1481
rect -1900 570 -1894 2593
rect 785 562 792 3203
rect 1152 3203 1202 3207
rect 4669 3180 7176 3186
rect 1123 3166 2074 3172
rect 2898 3105 3991 3106
rect 2701 3104 3991 3105
rect 2721 3094 3991 3104
rect 3998 3094 4000 3106
rect 2120 3062 5068 3073
rect 3683 3047 5153 3055
rect 976 2833 1015 2839
rect 4759 1418 5106 1426
rect 4759 1417 5121 1418
rect 2512 607 2516 769
rect 3096 607 3099 608
rect 2512 598 3099 607
rect 785 556 2236 562
rect 785 552 2183 556
rect 709 519 723 527
rect 730 519 788 527
rect -5371 472 -5367 477
rect -5113 473 -5110 478
rect -4606 235 -4598 440
rect -4146 426 -4105 427
rect -4146 416 -4130 426
rect -4110 416 -4105 426
rect -3807 422 -3795 429
rect -4146 -1131 -4105 416
rect -3821 -678 -3795 422
rect -3539 411 -3529 425
rect -3561 -515 -3529 411
rect -3301 398 -3261 403
rect -3274 -285 -3261 398
rect -69 203 -63 204
rect -69 194 14 203
rect 165 196 415 207
rect 702 203 709 519
rect 1112 426 1116 431
rect 2114 425 2115 430
rect 3096 430 3099 598
rect 5141 550 5153 3047
rect 7164 3002 7176 3180
rect 7164 1546 7176 2988
rect 7656 1655 7662 3387
rect 13000 3386 13117 3387
rect 13048 2487 13117 3386
rect 12740 2466 13117 2487
rect 13048 2424 13117 2466
rect 12796 2310 12800 2315
rect 11861 2249 12381 2253
rect 11902 2228 12381 2249
rect 8570 1644 10164 1653
rect 8122 1586 8124 1591
rect 8368 1587 8369 1592
rect 7708 1559 7709 1565
rect 7991 1560 8025 1564
rect 8235 1559 8246 1563
rect 7164 1539 7633 1546
rect 10146 866 10164 1644
rect 9890 857 10164 866
rect 10146 853 10164 857
rect 8488 766 8494 771
rect 8980 764 8981 769
rect 9921 763 10031 769
rect 9253 741 9259 750
rect 8980 724 8992 731
rect 8471 713 8472 720
rect 3060 424 3101 430
rect 846 339 1163 340
rect 846 326 1140 339
rect 846 324 1163 326
rect 1390 310 1397 416
rect 1592 334 8214 335
rect 1600 327 8214 334
rect 8241 327 8242 335
rect 1099 300 1101 306
rect 1108 300 1327 306
rect 1389 298 1398 310
rect 1555 300 7958 306
rect 841 285 875 290
rect 859 265 1313 270
rect 566 197 789 203
rect 940 195 1171 202
rect -180 49 -174 52
rect -69 50 -63 194
rect 209 135 212 140
rect 610 137 611 142
rect 984 134 985 139
rect 1356 125 1357 130
rect 844 104 862 106
rect 170 90 410 96
rect 571 94 574 98
rect 1390 98 1397 298
rect 7700 270 7703 274
rect 1570 265 7703 270
rect 7716 265 7751 274
rect 8471 240 8488 713
rect 1618 231 8491 240
rect 1606 228 8491 231
rect 7707 227 8491 228
rect 1214 96 1227 97
rect 571 91 784 94
rect 945 91 1140 94
rect 1135 85 1139 91
rect 1343 92 1397 98
rect 1135 82 1156 85
rect -180 43 -119 49
rect -180 -53 -174 43
rect -163 7 -145 13
rect -128 7 -113 13
rect -69 8 -27 14
rect 43 9 805 17
rect 431 -29 1175 -28
rect -128 -37 431 -33
rect 444 -37 1175 -29
rect 431 -38 1175 -37
rect -173 -60 -118 -53
rect -162 -96 -112 -90
rect -68 -95 -17 -89
rect -145 -153 -131 -96
rect -145 -168 844 -153
rect -131 -170 844 -168
rect 862 -169 1214 -153
rect 862 -170 1227 -169
rect 533 -285 539 -282
rect -3274 -294 539 -285
rect -3274 -297 -322 -294
rect -3274 -305 -1182 -297
rect 533 -374 539 -294
rect 8966 -304 8992 724
rect 513 -379 539 -374
rect 361 -399 370 -396
rect -3561 -557 2662 -515
rect 4802 -515 6925 -507
rect 2685 -551 8742 -515
rect 2685 -557 4810 -551
rect -3527 -559 4810 -557
rect 6920 -559 8742 -551
rect 9253 -671 9284 741
rect 9516 717 9527 725
rect 9542 717 9561 725
rect 9516 -512 9561 717
rect 9516 -556 9517 -512
rect 9516 -573 9561 -556
rect -3821 -680 -3733 -678
rect -3834 -750 2394 -680
rect 2417 -737 2418 -680
rect 2417 -738 2494 -737
rect 9253 -738 9277 -671
rect 2417 -750 9277 -738
rect -3834 -757 -3733 -750
rect -3834 -769 -3804 -757
rect -4108 -1186 -4105 -1131
<< m2contact >>
rect 11643 6740 11684 6751
rect 11573 6704 11601 6718
rect 12228 5413 12234 5427
rect 12278 5413 12283 5427
rect 8369 5245 8374 5254
rect 8634 5245 8667 5255
rect 1402 4513 1411 4521
rect 1431 4509 1454 4515
rect 3165 4017 3181 4023
rect 12381 3933 12387 3946
rect 12432 3933 12438 3947
rect 8124 3637 8132 3654
rect 12381 3637 12388 3654
rect -3241 2804 -3234 2809
rect -5346 2796 -5339 2801
rect -9788 2789 -9782 2794
rect -7479 2781 -7472 2786
rect -10370 2153 -10363 2178
rect -10798 1876 -10765 1906
rect -6598 1729 -6560 1763
rect -10797 1235 -10772 1281
rect -8893 1289 -8871 1324
rect -4476 1667 -4471 1674
rect -4476 1570 -4471 1579
rect -6598 1314 -6560 1356
rect -3989 589 -3984 595
rect -3686 591 -3681 598
rect -3419 587 -3414 595
rect -5243 505 -5238 510
rect -4985 506 -4980 511
rect -4733 508 -4726 513
rect -4476 507 -4471 512
rect -3989 505 -3984 510
rect -3686 508 -3681 513
rect -3419 505 -3414 510
rect 2701 3094 2721 3104
rect 969 2833 976 2839
rect 1015 2833 1021 2839
rect 1137 2833 1142 2839
rect 4730 1417 4759 1426
rect 5106 1418 5121 1426
rect 702 519 709 526
rect -4606 474 -4598 479
rect -3294 471 -3275 476
rect -4606 440 -4598 445
rect -3307 398 -3301 403
rect 983 458 988 463
rect 12507 2242 12513 2256
rect 8124 1586 8132 1591
rect 8369 1587 8374 1592
rect 8621 1583 8627 1588
rect 7657 1555 7666 1563
rect 7937 1556 7950 1564
rect 8182 1557 8195 1567
rect 8435 1553 8448 1563
rect 8563 1538 8575 1544
rect 7838 797 7845 802
rect 8100 798 8107 803
rect 8356 800 8361 805
rect 8611 799 8616 804
rect 8472 766 8488 771
rect 8966 764 8980 769
rect 9259 767 9284 773
rect 9527 764 9542 769
rect 10031 763 10041 769
rect 9259 741 9284 750
rect 8966 724 8980 731
rect 8472 713 8488 720
rect 985 134 991 139
rect 1357 125 1363 130
rect 30 105 43 114
rect 431 107 444 116
rect 62 99 85 107
rect 464 101 494 109
rect 805 104 818 110
rect 844 98 862 104
rect 1177 95 1190 104
rect 1214 89 1227 96
rect -145 7 -128 13
rect -27 8 -19 14
rect 30 9 43 17
rect 805 9 818 17
rect -145 -37 -128 -31
rect 431 -37 444 -29
rect 1175 -38 1190 -28
rect -181 -60 -173 -53
rect -17 -95 -11 -89
rect 844 -170 862 -153
rect 1214 -169 1227 -153
rect 265 -351 276 -344
rect 8965 -419 8992 -304
rect 9527 717 9542 725
<< metal2 >>
rect 11684 6740 11685 6749
rect 11573 6718 11601 6734
rect -3242 5924 -3233 5926
rect 11573 5924 11601 6704
rect -3242 5908 11601 5924
rect -3242 5350 -3233 5908
rect 11644 5865 11685 6740
rect 11644 5857 11686 5865
rect 8621 5846 11686 5857
rect -3242 5349 -3232 5350
rect -5346 3815 -5339 3816
rect -12654 3772 -5339 3815
rect -12654 3766 -12581 3772
rect -12687 -3560 -12581 3766
rect -7479 3639 -7472 3646
rect -12282 3509 -7472 3639
rect -12233 -2908 -12096 3509
rect -9788 3027 -9782 3055
rect -11482 3016 -9782 3027
rect -11489 278 -11432 3016
rect -9788 2794 -9782 3016
rect -7479 2786 -7472 3509
rect -5346 2801 -5339 3772
rect -3241 3621 -3232 5349
rect 8369 5254 8374 5255
rect 1402 4375 1411 4513
rect 657 4374 1411 4375
rect 653 4369 1411 4374
rect -3241 2809 -3237 3621
rect -10798 2178 -10762 2182
rect -10798 2153 -10370 2178
rect -10798 1906 -10762 2153
rect -10765 1876 -10762 1906
rect -6601 1763 -6557 1924
rect -6601 1729 -6598 1763
rect -6560 1729 -6557 1763
rect -4476 1674 -4471 1864
rect -3432 1626 -2330 1641
rect -8894 1289 -8893 1324
rect -4734 1355 -4725 1362
rect -6560 1315 -4725 1355
rect -10772 1235 -10771 1280
rect -10794 599 -10771 1235
rect -8894 894 -8872 1289
rect -8896 887 -4982 894
rect -10796 593 -5238 599
rect -5243 510 -5238 593
rect -4985 589 -4982 887
rect -4734 605 -4725 1315
rect -4985 511 -4981 589
rect -4733 513 -4726 605
rect -4476 512 -4471 1570
rect -3989 510 -3984 589
rect -3686 513 -3681 591
rect -3419 510 -3414 587
rect -4606 445 -4598 474
rect -3294 476 -3275 477
rect -3294 427 -3275 471
rect -2335 462 -2330 1626
rect -3203 427 -3165 429
rect -3294 426 -3165 427
rect -3293 422 -3165 426
rect -3203 389 -3165 422
rect -11489 276 -11425 278
rect -11482 -2376 -11425 276
rect -3204 -1356 -3111 389
rect -1805 299 -1796 1510
rect 653 356 657 4369
rect 1442 4225 1452 4509
rect 1442 4215 3190 4225
rect 3165 4023 3181 4215
rect 8124 3654 8128 3656
rect 702 2833 969 2839
rect 702 526 709 2833
rect 983 463 988 3264
rect 1036 3129 2749 3133
rect 1026 3101 2701 3104
rect 1037 3094 2701 3101
rect 1037 3093 2721 3094
rect 1021 2833 1137 2839
rect 2843 1426 2849 1429
rect 5474 1426 5497 1943
rect 8124 1591 8128 3637
rect 8369 1592 8374 5245
rect 8621 1588 8627 5846
rect 11644 5843 11686 5846
rect 12227 5413 12228 5427
rect 12227 5255 12234 5413
rect 8667 5245 12236 5255
rect 12278 5035 12283 5413
rect 14298 5035 14433 5048
rect 12275 5018 14433 5035
rect 12282 5017 14433 5018
rect 12387 3933 12388 3946
rect 12381 3654 12388 3933
rect 12432 3258 12436 3933
rect 13511 3258 13714 3318
rect 12432 3257 13714 3258
rect 12397 3249 13714 3257
rect 12397 3248 12433 3249
rect 12506 2256 12513 2257
rect 12506 2242 12507 2256
rect 2843 1417 4730 1426
rect 5121 1418 5496 1426
rect 5106 1417 5496 1418
rect 7657 1418 7666 1555
rect 2843 1415 4759 1417
rect 2843 944 2849 1415
rect 7657 1413 7845 1418
rect 2819 935 2826 939
rect 7838 802 7845 1413
rect 7943 1413 7947 1556
rect 8181 1557 8182 1567
rect 8100 1413 8107 1415
rect 7943 1404 8107 1413
rect 8100 803 8107 1404
rect 8181 1406 8195 1557
rect 8356 1406 8361 1409
rect 8181 1399 8361 1406
rect 8356 805 8361 1399
rect 8435 1398 8448 1553
rect 8575 1538 10041 1544
rect 8434 1390 8616 1398
rect 8611 804 8616 1390
rect 10030 1342 10041 1538
rect 8472 720 8488 766
rect 8966 731 8980 764
rect 10031 769 10041 1342
rect 9259 750 9284 767
rect 9527 725 9542 764
rect 653 351 802 356
rect -1805 295 617 299
rect 611 223 617 295
rect 985 139 992 351
rect 991 134 992 139
rect 7669 130 7677 690
rect 1363 125 7677 130
rect 30 17 43 105
rect -19 9 30 14
rect -19 7 43 9
rect -145 -31 -128 7
rect -181 -53 -173 -52
rect -181 -344 -173 -60
rect 71 -89 74 99
rect 431 -29 444 107
rect 470 -89 479 101
rect 805 17 818 104
rect -11 -95 487 -89
rect 844 -153 862 98
rect 1175 95 1177 104
rect 1175 -28 1190 95
rect 1214 -153 1227 89
rect -181 -351 265 -344
rect -181 -357 -173 -351
rect 8939 -419 8965 -304
rect 8992 -419 9007 -304
rect 8939 -570 9007 -419
rect 8940 -1084 9005 -570
rect 8940 -1108 9004 -1084
rect 2070 -1131 9004 -1108
rect 2115 -1178 9004 -1131
rect 2070 -1182 9004 -1178
rect 12506 -2376 12513 2242
rect -11482 -2462 12538 -2376
rect -11425 -2474 12538 -2462
rect 13511 -2511 13714 3249
rect 13511 -2908 13712 -2511
rect -12233 -3187 13712 -2908
rect -12105 -3219 13712 -3187
rect 14298 -3063 14433 5017
rect 14298 -3560 14422 -3063
rect -12687 -3691 14422 -3560
rect -12578 -3712 14422 -3691
<< m3contact >>
rect -5925 2271 -5911 2277
rect -6602 1924 -6557 1957
rect -4476 1864 -4471 1870
rect -1805 1510 -1796 1545
rect -2335 457 -2330 462
rect 3968 4021 3976 4029
rect 983 3264 993 3270
rect 1026 3129 1036 3139
rect 2749 3129 2754 3139
rect 1026 3093 1037 3101
rect 5474 1943 5497 1986
rect 611 218 617 223
rect 2070 -1178 2115 -1131
rect -3204 -1544 -3110 -1356
<< m123contact >>
rect 12288 6688 12305 6700
rect 1366 4498 1375 4503
rect -8063 2256 -8044 2263
rect -3823 2258 -3816 2267
rect -8893 1649 -8871 1680
rect -3203 565 -3197 570
rect -5386 472 -5381 477
rect -5129 473 -5113 478
rect -4864 475 -4854 480
rect -4130 472 -4110 477
rect -3827 475 -3808 480
rect -3560 472 -3541 477
rect -4130 416 -4110 426
rect -3828 422 -3807 429
rect -3198 459 -3192 465
rect -1900 565 -1894 570
rect -3562 411 -3539 426
rect -4606 225 -4598 235
rect -4146 -1186 -4108 -1131
rect 2017 3884 2037 3908
rect 785 3203 792 3208
rect 723 519 730 527
rect 1145 3201 1152 3209
rect 1202 3203 1208 3209
rect 1113 3166 1123 3172
rect 2074 3166 2083 3172
rect 3991 3094 3998 3106
rect 2112 3062 2120 3073
rect 5068 3062 5096 3073
rect 3668 3047 3683 3055
rect 7164 2988 7176 3002
rect 7837 1585 7845 1590
rect 12150 5419 12164 5434
rect 12512 5313 12532 5326
rect 12662 3833 12684 3846
rect 11861 2228 11902 2249
rect 12457 2242 12464 2256
rect 7709 1559 7725 1565
rect 7991 1553 8025 1560
rect 8228 1552 8246 1559
rect 8488 1555 8509 1561
rect 9098 797 9103 802
rect 9401 800 9414 805
rect 9669 797 9677 802
rect 9932 796 9939 801
rect 7703 764 7716 769
rect 7958 765 7981 770
rect 8214 767 8239 773
rect 9793 763 9817 768
rect 2236 556 2242 562
rect 5141 544 5153 550
rect 1240 459 1246 464
rect 1494 461 1500 466
rect 1749 460 1755 465
rect 2236 458 2242 463
rect 2540 461 2545 466
rect 2807 458 2812 463
rect 3071 457 3078 462
rect 775 426 780 432
rect 850 425 859 430
rect 1101 426 1108 431
rect 1353 428 1368 433
rect 1609 427 1628 432
rect 2096 425 2114 430
rect 2399 428 2418 433
rect 2666 425 2685 430
rect 2932 424 2951 429
rect 829 324 846 340
rect 832 285 841 290
rect 875 285 884 290
rect 840 265 859 270
rect 212 135 219 140
rect 611 137 617 142
rect 1140 326 1164 339
rect 1592 327 1600 334
rect 1101 300 1108 306
rect 1327 300 1338 306
rect 1542 300 1555 306
rect 1313 265 1328 270
rect 1557 265 1570 270
rect 1606 231 1618 240
rect 8214 326 8241 335
rect 7958 300 7982 306
rect 7703 265 7716 274
rect 13 90 21 96
rect -65 -26 -56 -19
rect -64 -128 -55 -122
rect 361 -396 370 -391
rect 322 -413 337 -401
rect 287 -461 304 -450
rect 2662 -557 2685 -513
rect 8742 -560 8811 -514
rect 9517 -556 9564 -512
rect 2394 -750 2417 -677
rect 12738 2142 12761 2155
<< metal3 >>
rect 15039 6709 15197 6834
rect 12288 6700 15197 6709
rect 12305 6688 15197 6700
rect 12131 5419 12150 5434
rect 3968 4698 3977 4705
rect 12131 4698 12164 5419
rect 15039 5331 15197 6688
rect 12512 5326 15197 5331
rect 12532 5313 15197 5326
rect 12512 5311 15197 5313
rect 3968 4684 12162 4698
rect 1366 3968 1375 4498
rect 3968 4083 3977 4684
rect 3968 4029 3976 4083
rect 1366 3958 2042 3968
rect 2017 3908 2037 3958
rect 15039 3850 15197 5311
rect 12662 3846 15197 3850
rect 12684 3833 15197 3846
rect 993 3264 1164 3267
rect 792 3203 1145 3207
rect 846 3173 851 3176
rect 846 3172 1123 3173
rect 846 3166 1113 3172
rect -8287 2263 -8267 2268
rect -6084 2266 -5925 2277
rect -4220 2267 -4214 2268
rect -8287 2256 -8063 2263
rect -8893 1950 -8864 1956
rect -8287 1950 -8267 2256
rect -6084 1958 -6065 2266
rect -4220 2258 -3823 2267
rect -6600 1957 -6063 1958
rect -8893 1930 -8258 1950
rect -8893 1680 -8864 1930
rect -6557 1924 -6063 1957
rect -4220 1870 -4214 2258
rect -4471 1864 -4212 1870
rect -8871 1649 -8864 1680
rect -3364 1510 -1805 1545
rect 846 1270 851 3166
rect 921 3133 931 3134
rect 921 3129 1026 3133
rect 2754 3129 3027 3133
rect 921 1404 931 3129
rect 5192 3125 5201 3128
rect 4033 3117 5201 3125
rect 1026 2062 1037 3093
rect 3071 3047 3668 3055
rect 1025 2061 1045 2062
rect 1554 2061 1564 2088
rect 1025 2055 1564 2061
rect 1045 2054 1564 2055
rect 921 1392 1500 1404
rect 846 1266 1246 1270
rect -3197 565 -1900 570
rect -1894 565 730 570
rect 723 527 730 565
rect -3828 480 -3807 481
rect -5386 273 -5381 472
rect -5129 290 -5113 473
rect -4864 333 -4854 475
rect -4130 426 -4110 472
rect -3828 475 -3827 480
rect -3808 475 -3807 480
rect -3828 429 -3807 475
rect -3562 472 -3560 477
rect -3541 472 -3539 477
rect -3562 426 -3539 472
rect 1240 464 1246 1266
rect -3192 459 -2335 462
rect -2330 459 754 462
rect 1494 466 1500 1392
rect 1554 798 1564 2054
rect 1749 798 1755 801
rect 1553 792 1755 798
rect 1749 465 1755 792
rect 5068 583 5096 3062
rect 2540 580 5096 583
rect 2236 463 2242 556
rect 751 432 754 459
rect 2540 466 2545 580
rect 2807 544 5141 550
rect 2807 463 2812 544
rect 3078 461 4886 462
rect 5192 461 5201 3117
rect 15039 3002 15197 3833
rect 7176 2988 15197 3002
rect 12456 2242 12457 2256
rect 11862 1989 11901 2228
rect 10922 1986 11249 1989
rect 5465 1943 5474 1986
rect 5497 1985 11249 1986
rect 11578 1985 11905 1989
rect 5497 1947 11905 1985
rect 5497 1943 10917 1947
rect 10922 1946 11905 1947
rect 11248 1942 11575 1946
rect 7841 1759 8677 1760
rect 12456 1759 12464 2242
rect 15039 2159 15197 2988
rect 12738 2155 15197 2159
rect 12761 2142 15197 2155
rect 12738 2140 15197 2142
rect 12738 2139 15039 2140
rect 7841 1755 12468 1759
rect 7841 1590 7845 1755
rect 8676 1753 12468 1755
rect 7702 1553 7726 1559
rect 7702 913 7709 1553
rect 7982 937 7991 1560
rect 8228 1102 8232 1552
rect 8476 1475 8508 1555
rect 8475 1468 9939 1475
rect 9931 1263 9939 1468
rect 9669 1102 9673 1109
rect 8228 1094 9673 1102
rect 7980 933 9406 937
rect 9339 932 9406 933
rect 9098 913 9103 914
rect 7702 910 9103 913
rect 9098 802 9103 910
rect 9401 805 9406 932
rect 9669 802 9673 1094
rect 9932 801 9939 1263
rect 7958 770 7981 771
rect 7703 769 7716 770
rect 3078 457 5199 461
rect 3071 456 5199 457
rect 751 426 775 432
rect 762 333 829 340
rect -4864 324 829 333
rect -4864 319 763 324
rect -5131 285 832 290
rect -5131 284 841 285
rect 850 273 859 425
rect 1101 306 1108 426
rect 1368 428 1372 433
rect 1353 339 1372 428
rect 1164 334 1372 339
rect 1609 392 1628 427
rect 1164 327 1592 334
rect 1164 326 1353 327
rect 1338 300 1542 306
rect 1101 290 1108 300
rect 884 287 1108 290
rect 884 285 1101 287
rect -5386 270 859 273
rect -5386 265 840 270
rect 1328 265 1557 270
rect -5386 264 850 265
rect 1609 254 1615 392
rect 1608 243 1616 254
rect -240 242 1618 243
rect -1008 240 1618 242
rect -1008 235 1606 240
rect -4598 231 1606 235
rect -4598 226 527 231
rect -4598 225 -4593 226
rect 611 142 617 218
rect 2096 202 2114 425
rect 2398 428 2399 433
rect 13 -19 21 90
rect -56 -26 21 -19
rect 13 -113 21 -26
rect 13 -122 22 -113
rect -55 -126 22 -122
rect -55 -128 13 -126
rect 6 -450 12 -128
rect 212 -401 216 135
rect 611 -53 617 137
rect 610 -205 617 -53
rect 237 -210 617 -205
rect 237 -212 505 -210
rect 610 -211 617 -210
rect 238 -392 245 -212
rect 238 -396 361 -392
rect 212 -413 322 -401
rect 6 -461 287 -450
rect 6 -479 12 -461
rect 2094 -550 2116 202
rect 2398 61 2418 428
rect 2658 430 2687 431
rect 2658 425 2666 430
rect 2685 425 2687 430
rect 2396 -311 2416 61
rect 2093 -551 2116 -550
rect -4146 -1131 -4081 -1129
rect 2093 -1131 2114 -551
rect 2394 -677 2416 -311
rect 2658 -499 2687 425
rect 2932 346 2951 424
rect 2931 104 2951 346
rect 7703 274 7716 764
rect 7958 306 7981 765
rect 8239 767 8240 773
rect 8214 335 8240 767
rect 9784 763 9793 768
rect 2664 -513 2683 -499
rect 2664 -568 2683 -557
rect 2394 -752 2416 -750
rect 2924 -904 2951 104
rect 8744 -510 8939 -509
rect 9008 -510 9559 -509
rect 8744 -512 9559 -510
rect 8744 -514 9517 -512
rect 8811 -556 9517 -514
rect 8811 -557 9559 -556
rect 8811 -559 8939 -557
rect 9008 -559 9559 -557
rect -4108 -1133 -4081 -1131
rect -3582 -1133 2070 -1132
rect -4108 -1177 2070 -1133
rect -4108 -1186 -3582 -1177
rect -4082 -1187 -3582 -1186
rect -3324 -1544 -3204 -1358
rect 2921 -1358 2956 -904
rect -3110 -1359 2965 -1358
rect 9784 -1359 9817 763
rect -3110 -1544 9819 -1359
rect -3324 -1547 9819 -1544
rect 2976 -1555 9819 -1547
use enable  enable_1
timestamp 1700021586
transform 1 0 -5274 0 1 473
box -177 -75 2126 105
use fourbitadder  fourbitadder_0
timestamp 1699884650
transform 1 0 -10308 0 1 1605
box -682 -95 8158 1279
use enable  enable_0
timestamp 1700021586
transform 1 0 952 0 1 426
box -177 -75 2126 105
use not  not_0
timestamp 1698904140
transform 1 0 -104 0 1 -16
box -15 -9 48 66
use not  not_1
timestamp 1698904140
transform 1 0 -103 0 1 -119
box -15 -9 48 66
use and  and_0
timestamp 1699601116
transform 1 0 15 0 1 83
box -14 7 194 122
use and  and_1
timestamp 1699601116
transform 1 0 416 0 1 85
box -14 7 194 122
use and  and_2
timestamp 1699601116
transform 1 0 790 0 1 82
box -14 7 194 122
use and  and_3
timestamp 1699601116
transform 1 0 1162 0 1 73
box -14 7 194 122
use tor  tor_0
timestamp 1699809212
transform 1 0 355 0 1 -410
box -90 -51 158 73
use comparator  comparator_0
timestamp 1701531022
transform 1 0 1105 0 1 3195
box -139 -2493 3703 970
use bitand  bitand_0
timestamp 1699892983
transform 1 0 7901 0 1 1553
box -276 -15 720 104
use enable  enable_2
timestamp 1700021586
transform 1 0 7813 0 1 765
box -177 -75 2126 105
use newor  newor_0
timestamp 1701531022
transform 1 0 12329 0 1 2140
box 0 -6 467 354
use and  and_4
timestamp 1699601116
transform 1 0 1386 0 1 4491
box -14 7 194 122
use newor  newor_1
timestamp 1701531022
transform 1 0 12252 0 1 3831
box 0 -6 467 354
use newor  newor_2
timestamp 1701531022
transform 1 0 12099 0 1 5311
box 0 -6 467 354
use tor  tor_1
timestamp 1699809212
transform 1 0 12150 0 1 6740
box -90 -51 158 73
<< labels >>
rlabel metal1 -56 198 -53 200 1 vdd
rlabel metal1 296 91 299 93 1 gnd
rlabel metal1 -155 9 -152 11 1 s0
rlabel metal1 -157 -94 -154 -92 1 s1
rlabel metal1 614 139 615 140 1 d1
rlabel m2contact 988 136 989 137 1 d2
rlabel m2contact 1360 127 1361 128 7 d3
rlabel metal1 1581 4545 1582 4546 1 equal
rlabel metal2 2822 936 2823 937 1 big
rlabel m2contact -9783 2791 -9782 2792 1 sum0
rlabel m2contact -7474 2783 -7473 2784 1 sum1
rlabel m2contact -5341 2798 -5340 2799 1 sum2
rlabel metal1 -2187 2559 -2186 2560 1 sum4
rlabel m2contact 8372 1589 8373 1590 1 k2
rlabel metal1 7843 1587 7844 1588 1 k0
rlabel m2contact 8625 1585 8626 1586 1 k3
rlabel m2contact -3239 2806 -3238 2807 1 sum3
rlabel m2contact 8126 1588 8127 1589 1 k1
rlabel m3contact 3972 4026 3973 4027 1 small
rlabel metal1 12798 2312 12799 2313 1 final0
rlabel metal1 12721 4003 12722 4004 1 final1
rlabel metal1 12568 5483 12569 5484 1 final2
rlabel metal1 12310 6773 12311 6774 1 final3
rlabel m123contact -5384 473 -5383 474 1 aa0
rlabel m123contact -5119 474 -5118 475 1 aa1
rlabel m123contact -4858 476 -4857 477 1 aa2
rlabel m2contact -4602 475 -4601 476 1 aa3
rlabel m123contact -4118 474 -4117 475 1 bb0
rlabel m123contact -3816 477 -3815 478 1 bb1
rlabel m123contact -3544 473 -3543 474 1 bb2
rlabel m2contact -3280 473 -3279 474 1 bb3
rlabel metal1 3016 4025 3017 4026 1 eq1
<< end >>
