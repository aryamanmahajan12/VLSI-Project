* SPICE3 file created from and.ext - technology: scmos

.include TSMC_180nm.txt

.option scale=0.09u


.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd vdd gnd 'SUPPLY'



Vinb b gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)

Vina a gnd PULSE(0 1.8 0ns 100ps 100ps 30ns 50ns)





.option scale=0.09u

M1000 out not_0/in vdd not_0/w_n15_38# CMOSP w=7 l=4
+  ad=70 pd=34 as=733 ps=188
M1001 out not_0/in gnd Gnd CMOSN w=6 l=4
+  ad=60 pd=32 as=313 ps=100
M1002 not_0/in a vdd nand_0/w_n44_54# CMOSP w=13 l=9
+  ad=390 pd=86 as=0 ps=0
M1003 not_0/in b nand_0/a_n8_22# Gnd CMOSN w=11 l=3
+  ad=187 pd=56 as=330 ps=82
M1004 vdd b not_0/in nand_0/w_n44_54# CMOSP w=13 l=3
+  ad=0 pd=0 as=0 ps=0
M1005 nand_0/a_n8_22# a gnd Gnd CMOSN w=11 l=9
+  ad=0 pd=0 as=0 ps=0
C0 not_0/w_n15_38# vdd 0.09fF
C1 b nand_0/w_n44_54# 0.14fF
C2 out vdd 0.03fF
C3 not_0/w_n15_38# not_0/in 0.11fF
C4 nand_0/w_n44_54# a 0.28fF
C5 b not_0/in 0.10fF
C6 out not_0/w_n15_38# 0.04fF
C7 vdd nand_0/w_n44_54# 0.13fF
C8 not_0/in nand_0/w_n44_54# 0.06fF
C9 gnd Gnd 1.01fF
C10 not_0/in Gnd 0.82fF
C11 b Gnd 0.28fF
C12 a Gnd 0.53fF
C13 nand_0/w_n44_54# Gnd 3.07fF
C14 out Gnd 0.22fF
C15 not_0/w_n15_38# Gnd 1.29fF





.tran 1n 800n

.control

run
set color0 = rgb:f/f/e
set color1 = black

plot v(a) v(b)+4 v(out)+8

.end
.endc