magic
tech scmos
timestamp 1699876194
<< metal1 >>
rect 2742 696 3067 706
rect 2812 646 2825 651
rect 3061 628 3068 696
rect 3590 628 3609 629
rect 3212 618 3635 628
rect 3590 617 3635 618
rect 2208 270 2220 568
rect 3256 558 3534 564
rect 2272 437 2284 555
rect 3105 522 3106 530
rect 3038 514 3056 517
rect 2598 484 2628 494
rect 3026 508 3056 514
rect 3026 484 3038 508
rect 2598 461 3040 484
rect 2598 458 2628 461
rect 2780 437 2798 438
rect 2271 436 2798 437
rect 2271 404 2768 436
rect 2780 217 2798 404
rect 2194 -61 2218 136
rect 2256 4 2263 121
rect 2615 39 2633 60
rect 2913 39 2923 461
rect 3206 327 3216 513
rect 3521 377 3534 558
rect 3622 434 3634 617
rect 3863 435 3929 441
rect 3865 399 3881 404
rect 3709 379 3722 386
rect 3521 367 3698 377
rect 3534 365 3698 367
rect 3206 319 3639 327
rect 3206 308 3216 319
rect 3900 160 3924 435
rect 3232 138 3924 160
rect 3121 41 3122 49
rect 3152 41 3155 49
rect 2615 38 2923 39
rect 2615 31 3077 38
rect 2615 29 2923 31
rect 2615 12 2633 29
rect 2913 24 2923 29
rect 2256 -12 3098 4
rect 3111 -12 3112 4
rect 2256 -13 2263 -12
rect 3718 -61 3749 138
rect 3900 137 3924 138
rect 2194 -86 3762 -61
rect 2194 -88 2218 -86
<< m2contact >>
rect 3077 528 3090 539
rect 2598 494 2628 509
rect 2768 404 2798 436
rect 2615 60 2633 75
rect 3701 379 3709 386
rect 3268 77 3277 82
rect 3098 47 3111 55
rect 3098 -12 3111 4
<< metal2 >>
rect 3074 528 3077 539
rect 3090 528 3092 539
rect 3074 437 3092 528
rect 2769 436 3089 437
rect 2798 404 3089 436
rect 2769 403 3089 404
rect 3598 386 3616 389
rect 3598 379 3701 386
rect 3598 87 3616 379
rect 3268 82 3628 87
rect 3277 77 3628 82
rect 3098 4 3111 47
<< m123contact >>
rect 2309 571 2319 576
rect 3106 522 3140 530
rect 2305 137 2319 142
rect 3122 41 3152 49
<< metal3 >>
rect 2309 388 2319 571
rect 3106 388 3140 522
rect 2309 365 3124 388
rect 2318 361 3124 365
rect 2305 -20 2319 137
rect 3122 -20 3152 41
rect 2305 -32 3151 -20
use tor  tor_1
timestamp 1699809212
transform 1 0 3707 0 1 368
box -90 -51 158 73
use and  and_1
timestamp 1699601116
transform 1 0 3062 0 1 506
box -14 7 194 122
use and  and_0
timestamp 1699601116
transform 1 0 3083 0 1 25
box -14 7 194 122
use xor  xor_1
timestamp 1699082409
transform 1 0 2227 0 1 602
box -18 -108 585 124
use xor  xor_0
timestamp 1699082409
transform 1 0 2225 0 1 168
box -18 -108 585 124
<< labels >>
rlabel metal1 2210 326 2214 328 1 vdd
rlabel metal1 2764 33 2768 35 1 gnd
rlabel metal1 2266 -8 2270 -6 1 a
rlabel metal3 2311 26 2315 28 1 b
rlabel metal3 2455 369 2459 371 1 c
rlabel metal1 2820 647 2822 648 1 s
rlabel metal1 3873 400 3875 401 1 carry
<< end >>
