magic
tech scmos
timestamp 1699884650
<< metal1 >>
rect 749 1248 1625 1249
rect 2164 1248 2216 1250
rect -278 1211 -108 1248
rect 749 1234 2216 1248
rect 749 1233 2163 1234
rect 1626 1232 2163 1233
rect 3057 1226 4337 1236
rect 5196 1222 6438 1233
rect -261 1210 -201 1211
rect -261 203 -202 1210
rect 7054 1199 7066 1204
rect 4953 1191 4964 1196
rect 507 1184 522 1189
rect 2815 1176 2831 1181
rect 8110 952 8118 957
rect -56 686 -48 695
rect 4390 694 4399 704
rect 6491 700 6497 708
rect 2252 671 2265 682
rect 2727 236 4325 241
rect 4861 238 6454 248
rect 2727 229 4328 236
rect 4883 231 6454 238
rect 2725 220 4328 229
rect -261 196 -130 203
rect 402 198 2192 214
rect -261 192 -131 196
rect -202 189 -131 192
rect 4383 120 4389 126
rect 2247 106 2253 112
rect 6478 114 6484 120
rect -76 84 -70 90
<< metal2 >>
rect -682 1026 -91 1062
rect -609 642 -558 1026
rect -609 624 -92 642
rect 4043 627 4131 629
rect -609 20 -558 624
rect 1848 619 1904 620
rect 1848 572 2215 619
rect 4043 592 4353 627
rect 6210 624 6455 632
rect 6166 596 6455 624
rect -609 7 -112 20
rect -609 6 -558 7
rect 322 6 1672 7
rect 1848 6 1904 572
rect 4043 49 4131 592
rect 6166 49 6209 596
rect 2646 48 4347 49
rect 2122 6 2210 29
rect 2645 17 4347 48
rect 4781 18 6441 49
rect 322 -6 2210 6
rect 1672 -7 2210 -6
<< m123contact >>
rect 5994 943 6009 949
rect 1551 937 1563 942
rect 3859 929 3871 934
rect 446 146 472 151
rect -29 71 -15 76
rect 2769 169 2794 174
rect 2288 94 2299 99
rect 4906 186 4927 191
rect 4431 111 4438 116
rect 7001 173 7025 178
rect 6524 98 6539 103
<< metal3 >>
rect 6153 1023 6538 1024
rect -313 1007 -9 1013
rect 4145 1009 4437 1012
rect -387 968 -9 1007
rect 2015 976 2299 1004
rect 4128 997 4437 1009
rect 6139 1004 6538 1023
rect -387 701 -315 968
rect 2015 945 2031 976
rect 1551 942 2031 945
rect 1563 937 2031 942
rect 4128 934 4145 997
rect 6139 949 6153 1004
rect 6009 943 6161 949
rect 3871 929 4145 934
rect -387 651 -316 701
rect -387 625 -317 651
rect -387 -57 -316 625
rect 446 151 472 506
rect 2769 174 2794 498
rect 4906 191 4927 513
rect 7001 178 7025 521
rect 2299 94 2300 99
rect -29 -57 -15 71
rect -417 -58 -15 -57
rect 2288 -58 2300 94
rect -417 -61 3962 -58
rect 4431 -61 4438 111
rect -417 -62 4956 -61
rect 6524 -62 6539 98
rect -417 -89 6944 -62
rect -29 -90 6944 -89
rect -14 -91 6944 -90
rect 3962 -94 6944 -91
rect 4956 -95 6944 -94
use xor  xor_0
timestamp 1699082409
transform 1 0 -113 0 1 102
box -18 -108 585 124
use fulladder  fulladder_0
timestamp 1699876194
transform 1 0 -2318 0 1 538
box 2194 -88 3929 726
use xor  xor_1
timestamp 1699082409
transform 1 0 2210 0 1 125
box -18 -108 585 124
use fulladder  fulladder_1
timestamp 1699876194
transform 1 0 -10 0 1 530
box 2194 -88 3929 726
use xor  xor_2
timestamp 1699082409
transform 1 0 4346 0 1 142
box -18 -108 585 124
use fulladder  fulladder_2
timestamp 1699876194
transform 1 0 2128 0 1 545
box 2194 -88 3929 726
use xor  xor_3
timestamp 1699082409
transform 1 0 6441 0 1 129
box -18 -108 585 124
use fulladder  fulladder_3
timestamp 1699876194
transform 1 0 4229 0 1 553
box 2194 -88 3929 726
<< labels >>
rlabel metal3 -372 227 -362 252 1 m
rlabel metal2 -593 284 -585 298 1 gnd
rlabel metal1 -241 300 -233 314 1 vdd
rlabel metal1 -75 86 -73 87 1 b0
rlabel metal1 2249 109 2251 110 1 b1
rlabel metal1 4385 123 4387 124 1 b2
rlabel metal1 6481 116 6483 117 1 b3
rlabel metal1 -54 689 -52 691 1 a0
rlabel metal1 2257 675 2260 677 1 a1
rlabel metal1 4392 697 4393 699 1 a2
rlabel metal1 6492 703 6494 704 1 a3
rlabel metal1 516 1185 519 1187 1 s0
rlabel metal1 2820 1178 2822 1179 1 s1
rlabel metal1 4959 1192 4960 1193 1 s2
rlabel metal1 7059 1201 7061 1202 1 s3
rlabel metal1 8114 954 8115 955 1 s4
<< end >>
